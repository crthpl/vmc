module packets
