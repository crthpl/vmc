module packets

pub type Packet = Handshake | Ping | Request
