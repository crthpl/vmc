module packets

pub struct Packeter {
pub:
	server bool
pub mut:
	version int = -1
}
